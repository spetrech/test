module  top();
endmodule
